-------------------------------------------------------------
--
-- Lab 01
--
-- Written By Jim Lynch
-- 01.10.2023
--
-------------------------------------------------------------